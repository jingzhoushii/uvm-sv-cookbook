// ============================================================================
// Testbench: tb_data_types
// 功能: 验证 SystemVerilog 数据类型的特性和用法
// ============================================================================
`timescale 1ns/1ps

module tb_data_types;
    // ------------------------------------------------------------------------
    // 时钟和复位信号
    // ------------------------------------------------------------------------
    reg  clk;           // 系统时钟，周期 10ns
    reg  rst_n;         // 低电平复位信号，异步复位
    
    // ------------------------------------------------------------------------
    // ALU 接口信号
    // ------------------------------------------------------------------------
    reg  [31:0] a;         // 操作数 A
    reg  [31:0] b;         // 操作数 B
    reg  [3:0]  opcode;    // 操作码：定义 ALU 执行的操作类型
    wire [31:0] result;    // 计算结果输出
    
    // ------------------------------------------------------------------------
    // 实例化被测设计 (DUT)
    // ------------------------------------------------------------------------
    simple_alu dut (
        .clk(clk),         // 时钟输入
        .rst_n(rst_n),     // 复位输入（低有效）
        .a(a),             // 操作数 A
        .b(b),             // 操作数 B
        .opcode(opcode),   // 操作码
        .result(result)     // 结果输出
    );
    
    // ------------------------------------------------------------------------
    // 时钟生成器
    // 周期: 10ns (频率: 100MHz)
    // ------------------------------------------------------------------------
    initial begin
        clk = 0;
        forever #5 clk = ~clk;  // 每 5ns 翻转一次
    end
    
    // ------------------------------------------------------------------------
    // 复位和测试激励序列
    // ------------------------------------------------------------------------
    initial begin
        // 1. 复位阶段
        rst_n = 0;          // 断言复位
        #10 rst_n = 1;      // 10ns 后释放复位
        
        // 2. 测试用例 1: 加法 (opcode=0)
        a = 10;             // 设置操作数 A
        b = 5;              // 设置操作数 B
        opcode = 0;         // 加法操作
        #10;                // 等待一个时钟周期
        
        // 3. 测试用例 2: 减法 (opcode=1)
        opcode = 1;         // 减法操作
        #10;
        
        // 4. 测试用例 3: 乘法 (opcode=2)
        opcode = 2;         // 乘法操作
        #30;                // 等待 30ns 观察结果
        
        // 5. 结束仿真
        $finish;
    end
    
    // ------------------------------------------------------------------------
    // 波形记录
    // 用于 EDA 工具（如 GTKwave, Verdi）查看信号波形
    // ------------------------------------------------------------------------
    initial begin
        $dumpfile("dump.vcd");           // 指定波形文件
        $dumpvars(0, tb_data_types);     // 记录模块中所有信号
    end
    
endmodule
