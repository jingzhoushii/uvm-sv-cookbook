// ============================================================================
// SystemVerilog OOP 示例 - 格式化版本
// ============================================================================
// 本文件展示 SystemVerilog 面向对象编程的核心概念
// ============================================================================

`timescale 1ns/1ps

// ============================================================================
// 基类：base
// 功能：演示基本的类定义、构造函数和虚函数
// ============================================================================
class base;
    int x;  // 成员变量
    
    // ------------------------------------------------------------------------
    // 构造函数
    // ------------------------------------------------------------------------
    function new(int v);
        x = v;  // 初始化成员变量
    endfunction
    
    // ------------------------------------------------------------------------
    // 虚函数：支持多态
    // ------------------------------------------------------------------------
    virtual function void disp();
        $display("base: x=%0d", x);
    endfunction
endclass

// ============================================================================
// 派生类：derived
// 功能：演示继承和方法覆盖
// ============================================================================
class derived extends base;
    int y;  // 新增成员变量
    
    // ------------------------------------------------------------------------
    // 构造函数：调用父类构造函数
    // ------------------------------------------------------------------------
    function new(int a, int b);
        super.new(a);  // 调用父类构造函数
        y = b;         // 初始化新变量
    endfunction
    
    // ------------------------------------------------------------------------
    // 覆盖父类的 disp() 方法
    // ------------------------------------------------------------------------
    virtual function void disp();
        $display("derived: x=%0d y=%0d", x, y);
    endfunction
endclass

// ============================================================================
// 测试模块
// 功能：演示多态和类型转换
// ============================================================================
module tb_oop;
    initial begin
        // 1. 创建基类和派生类对象
        base     b;       // 基类句柄
        derived  d;       // 派生类对象
        
        b = new(10);          // 创建基类对象
        d = new(20, 30);      // 创建派生类对象
        
        // 2. 调用方法
        b.disp();             // 调用 base::disp() → "base: x=10"
        d.disp();             // 调用 derived::disp() → "derived: x=20 y=30"
        
        // 3. 多态演示：基类句柄指向派生类对象
        b = d;                // 父类句柄指向子类对象
        
        // 4. 类型转换：安全地将基类句柄转回派生类
        $cast(d, b);          // 运行时类型检查
        
        // 5. 再次调用：仍然是派生类的方法
        d.disp();             // "derived: x=20 y=30"
        
        // 6. 结束仿真
        #100;
        $finish;
    end
    
    // ------------------------------------------------------------------------
    // 波形记录
    // ------------------------------------------------------------------------
    initial begin
        $dumpfile("dump.vcd");
        $dumpvars(0, tb_oop);
    end
endmodule
