// ============================================================================
// SystemVerilog Interfaces 示例 - 格式化版本
// ============================================================================
// 本文件展示 SystemVerilog 接口的定义和使用
// ============================================================================

`timescale 1ns/1ps

// ============================================================================
// 总线接口：bus_if
// 功能：封装总线信号和协议操作
// 信号：addr, data, rw, valid, ready
// ============================================================================
interface bus_if (input bit clk);
    // ------------------------------------------------------------------------
    // 信号声明
    // ------------------------------------------------------------------------
    logic [31:0] addr;    // 地址总线
    logic [31:0] data;    // 数据总线
    logic         rw;      // 读写控制：1=写，0=读
    logic         valid;   // 有效信号
    logic         ready;   // 就绪信号（从设备产生）
    
    // ------------------------------------------------------------------------
    // modport：定义信号方向
    // ------------------------------------------------------------------------
    modport master (
        output addr,        // 主设备输出地址
        output data,        // 主设备输出数据
        output rw,          // 主设备输出读写控制
        output valid,       // 主设备输出有效信号
        input  ready       // 主设备输入就绪信号
    );
    
    modport slave (
        input  addr,        // 从设备输入地址
        input  data,        // 从设备输入数据
        input  rw,          // 从设备输入读写控制
        input  valid,       // 从设备输入有效信号
        output ready        // 从设备输出就绪信号
    );
    
    // ------------------------------------------------------------------------
    // 任务：主设备写操作
    // 协议：发起传输 → 等待就绪 → 完成
    // ------------------------------------------------------------------------
    task master_write(
        input [31:0] a,  // 地址参数
        input [31:0] d   // 数据参数
    );
        // 1. 放置地址和数据
        addr  = a;
        data  = d;
        rw    = 1;       // 写操作
        valid = 1;       // 断言有效
        
        // 2. 等待时钟上升沿采样
        @(posedge clk);
        
        // 3. 等待从设备就绪
        while (!ready) begin
            @(posedge clk);
        end
        
        // 4. 结束传输
        valid = 0;
    endtask
endinterface

// ============================================================================
// 测试模块
// 功能：演示接口的使用
// ============================================================================
module tb_if;
    bit clk;                    // 系统时钟
    bus_if ifc(clk);           // 接口实例
    
    // ------------------------------------------------------------------------
    // 时钟生成器
    // ------------------------------------------------------------------------
    initial begin
        clk = 0;
        forever #5 clk = ~clk;  // 周期：10ns
    end
    
    // ------------------------------------------------------------------------
    // 测试序列
    // ------------------------------------------------------------------------
    initial begin
        // 等待复位稳定
        #10;
        
        // 执行一次写操作
        ifc.master_write(32'h1000, 32'hABCD);
        
        // 仿真结束
        #100;
        $finish;
    end
    
    // ------------------------------------------------------------------------
    // 波形记录
    // ------------------------------------------------------------------------
    initial begin
        $dumpfile("dump.vcd");
        $dumpvars(0, tb_if);
    end
endmodule
