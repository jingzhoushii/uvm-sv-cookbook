// ============================================================================
// SystemVerilog Randomization 示例 - 格式化版本
// ============================================================================
// 本文件展示 SystemVerilog 随机化和约束的使用
// ============================================================================

`timescale 1ns/1ps

// ============================================================================
// Transaction 类
// 功能：带约束的随机事务生成
// ============================================================================
class tx;
    // ------------------------------------------------------------------------
    // 随机变量
    // ------------------------------------------------------------------------
    rand bit [7:0] d;     // 数据：0-255
    rand bit [3:0] len;  // 长度：0-15
    
    // ------------------------------------------------------------------------
    // 约束 c1：范围约束
    // 功能：限制 d 和 len 的取值范围
    // ------------------------------------------------------------------------
    constraint c1 {
        d inside {[10:100]};    // 数据在 10-100 之间
        len inside {[1:10]};    // 长度在 1-10 之间
    }
    
    // ------------------------------------------------------------------------
    // 约束 c2：条件约束（Implication）
    // 功能：当 d>50 时，len<5
    // 语法：条件 -> 结果
    // ------------------------------------------------------------------------
    constraint c2 {
        d > 50 -> len < 5;
    }
    
    // ------------------------------------------------------------------------
    // 约束 c3：分布约束
    // 功能：控制各取值的概率分布
    // 语法：值 dist {权重}
    // ------------------------------------------------------------------------
    constraint c3 {
        len dist {
            0 :/ 10,   // len=0 的权重：10
            1 :/ 30,   // len=1 的权重：30
            2 :/ 60    // len=2 的权重：60
        };
    }
endclass

// ============================================================================
// 测试模块
// 功能：演示随机化调用
// ============================================================================
module tb_rnd;
    initial begin
        tx t;
        
        $display("========================================");
        $display("  SystemVerilog Randomization Demo");
        $display("========================================");
        
        t = new();
        
        // 生成 5 个随机事务
        repeat (5) begin
            // 随机化并检查结果
            if (t.randomize()) begin
                $display("d=%0d  len=%0d", t.d, t.len);
            end else begin
                $display("ERROR: Randomization failed!");
            end
            
            #10;  // 间隔 10ns
        end
        
        $display("\nRandomization test Complete!");
        #100;
        $finish;
    end
    
    // ------------------------------------------------------------------------
    // 波形记录
    // ------------------------------------------------------------------------
    initial begin
        $dumpfile("dump.vcd");
        $dumpvars(0, tb_rnd);
    end
endmodule
