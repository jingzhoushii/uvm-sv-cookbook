// ============================================================================
// Testbench: tb_interfaces
// 功能: 验证 SystemVerilog Interface 的使用方法
// 知识点: modport, interface, clocking block
// ============================================================================
`timescale 1ns/1ps

module tb_interfaces;
    // ------------------------------------------------------------------------
    // 接口信号
    // ------------------------------------------------------------------------
    bit  clk;              // 系统时钟，周期 10ns
    bit  rst_n;           // 低电平复位信号
    
    // ------------------------------------------------------------------------
    // 实例化总线接口
    // bus_if 包含: addr, data, rw, valid, ready 等信号
    // ------------------------------------------------------------------------
    bus_if ifc (clk, rst_n);  // 接口实例，连接到时钟和复位
    
    // ------------------------------------------------------------------------
    // 驱动器 (Driver)：产生测试激励
    // ------------------------------------------------------------------------
    initial begin
        // 1. 初始化
        clk = 0;
        forever #5 clk = ~clk;  // 时钟生成：100MHz
    end
    
    // ------------------------------------------------------------------------
    // 复位和测试序列
    // ------------------------------------------------------------------------
    initial begin
        // 复位阶段
        rst_n = 0;
        #10 rst_n = 1;
        
        // 发送 5 个写事务
        repeat (5) begin
            // 产生随机地址和数据
            ifc.addr = $random & 32'h00FF;  // 限制地址范围
            ifc.wdata = $random;            // 随机写数据
            ifc.valid = 1'b1;                // 断言有效信号
            
            // 等待时钟上升沿采样
            @(posedge clk);
            #1;  // 延迟 1ns 确保稳定
            
            // 打印事务信息
            $display("addr=0x%0h wdata=0x%0h valid=%0d",
                     ifc.addr, ifc.wdata, ifc.valid);
            
            // 等待总线就绪（如果有 ready 信号）
            // while (!ifc.ready) @(posedge clk);
        end
        
        // 测试完成
        $display("Interface Demo Complete!");
        $finish;
    end
    
    // ------------------------------------------------------------------------
    // 波形记录
    // ------------------------------------------------------------------------
    initial begin
        $dumpfile("dump.vcd");
        $dumpvars(0, tb_interfaces);
    end
    
endmodule
